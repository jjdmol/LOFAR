-- megafunction wizard: %FFT-IFFT v1.3.0%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: aukfft_core 

-- ============================================================
-- File Name: myfftcore.vhd
-- Megafunction Name(s):
-- 			aukfft_core
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
-- ************************************************************


--Copyright (C) 1991-2002 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY myfftcore IS
	PORT
	(
		sysclk			: IN STD_LOGIC ;
		reset			: IN STD_LOGIC ;
		go				: IN STD_LOGIC ;
		realdatain		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
		imagdatain		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
		realtwid		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
		imagtwid		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
		realdataout		: OUT STD_LOGIC_VECTOR (16 DOWNTO 1);
		imagdataout		: OUT STD_LOGIC_VECTOR (16 DOWNTO 1);
		readaddress		: OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		writeaddress	: OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		twidaddress		: OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		exponent		: OUT STD_LOGIC_VECTOR (5 DOWNTO 1);
		done			: OUT STD_LOGIC ;
		writeenable		: OUT STD_LOGIC ;
		direction		: OUT STD_LOGIC 
	);
END myfftcore;

ARCHITECTURE SYN OF myfftcore IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (8 DOWNTO 1);
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (16 DOWNTO 1);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (5 DOWNTO 1);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (8 DOWNTO 1);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (8 DOWNTO 1);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (16 DOWNTO 1);

	COMPONENT aukfft_core
	GENERIC (
		floatwidth			: NATURAL;
		datawidth			: NATURAL;
		twiddlewidth		: NATURAL;
		points				: NATURAL;
		stratix				: NATURAL;
		backward_compatible	: NATURAL;
		transform			: STRING;
		interface			: STRING
	);
	PORT (
			realdatain		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
			direction		: OUT STD_LOGIC ;
			done			: OUT STD_LOGIC ;
			writeaddress	: OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
			writeenable		: OUT STD_LOGIC ;
			imagtwid		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
			sysclk			: IN STD_LOGIC ;
			realtwid		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
			reset			: IN STD_LOGIC ;
			realdataout		: OUT STD_LOGIC_VECTOR (16 DOWNTO 1);
			go				: IN STD_LOGIC ;
			imagdatain		: IN STD_LOGIC_VECTOR (16 DOWNTO 1);
			exponent		: OUT STD_LOGIC_VECTOR (5 DOWNTO 1);
			twidaddress		: OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
			readaddress		: OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
			imagdataout		: OUT STD_LOGIC_VECTOR (16 DOWNTO 1)
	);
	END COMPONENT;

BEGIN
	direction    			<= sub_wire0;
	done    				<= sub_wire1;
	writeaddress    		<= sub_wire2(8 DOWNTO 1);
	writeenable    			<= sub_wire3;
	realdataout    			<= sub_wire4(16 DOWNTO 1);
	exponent    			<= sub_wire5(5 DOWNTO 1);
	twidaddress   	 		<= sub_wire6(8 DOWNTO 1);
	readaddress    			<= sub_wire7(8 DOWNTO 1);
	imagdataout    			<= sub_wire8(16 DOWNTO 1);

	aukfft_core_component : aukfft_core
	GENERIC MAP (
		floatwidth 			=> 4,
		datawidth 			=> 16,
		twiddlewidth 		=> 16,
		points 				=> 256,
		stratix 			=> 0,
		backward_compatible => 0,
		transform 			=> "fft",
		interface 			=> "internal"
	)
	PORT MAP (
		realdatain 			=> realdatain,
		imagtwid 			=> imagtwid,
		sysclk 				=> sysclk,
		realtwid 			=> realtwid,
		reset 				=> reset,
		go 					=> go,
		imagdatain 			=> imagdatain,
		direction 			=> sub_wire0,
		done 				=> sub_wire1,
		writeaddress 		=> sub_wire2,
		writeenable 		=> sub_wire3,
		realdataout 		=> sub_wire4,
		exponent 			=> sub_wire5,
		twidaddress 		=> sub_wire6,
		readaddress 		=> sub_wire7,
		imagdataout 		=> sub_wire8
	);

END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: DATAWIDTH NUMERIC 16
-- Retrieval info: PRIVATE: TWIDDLEWIDTH NUMERIC 16
-- Retrieval info: PRIVATE: POINTS NUMERIC 256
-- Retrieval info: PRIVATE: POINTSLOG2 NUMERIC 8
-- Retrieval info: PRIVATE: FLOATWIDTH NUMERIC 4
-- Retrieval info: PRIVATE: INTERNALMEM NUMERIC 1
-- Retrieval info: PRIVATE: FFT NUMERIC 1
-- Retrieval info: PRIVATE: STRATIX NUMERIC 0
-- Retrieval info: PRIVATE: BACKWARD_COMPATIBLE NUMERIC 0
-- Retrieval info: CONSTANT: floatwidth NUMERIC 4
-- Retrieval info: CONSTANT: datawidth NUMERIC 16
-- Retrieval info: CONSTANT: twiddlewidth NUMERIC 16
-- Retrieval info: CONSTANT: points NUMERIC 256
-- Retrieval info: CONSTANT: stratix NUMERIC 0
-- Retrieval info: CONSTANT: backward_compatible NUMERIC 0
-- Retrieval info: CONSTANT: transform STRING fft
-- Retrieval info: CONSTANT: interface STRING internal
-- Retrieval info: USED_PORT: sysclk 0 0 0 0 INPUT NODEFVAL sysclk
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL reset
-- Retrieval info: USED_PORT: go 0 0 0 0 INPUT NODEFVAL go
-- Retrieval info: USED_PORT: realdatain 0 0 16 1 INPUT NODEFVAL realdatain[16..1]
-- Retrieval info: USED_PORT: imagdatain 0 0 16 1 INPUT NODEFVAL imagdatain[16..1]
-- Retrieval info: USED_PORT: realtwid 0 0 16 1 INPUT NODEFVAL realtwid[16..1]
-- Retrieval info: USED_PORT: imagtwid 0 0 16 1 INPUT NODEFVAL imagtwid[16..1]
-- Retrieval info: USED_PORT: realdataout 0 0 16 1 OUTPUT NODEFVAL realdataout[16..1]
-- Retrieval info: USED_PORT: imagdataout 0 0 16 1 OUTPUT NODEFVAL imagdataout[16..1]
-- Retrieval info: USED_PORT: readaddress 0 0 8 1 OUTPUT NODEFVAL readaddress[8..1]
-- Retrieval info: USED_PORT: writeaddress 0 0 8 1 OUTPUT NODEFVAL writeaddress[8..1]
-- Retrieval info: USED_PORT: twidaddress 0 0 8 1 OUTPUT NODEFVAL twidaddress[8..1]
-- Retrieval info: USED_PORT: exponent 0 0 5 1 OUTPUT NODEFVAL exponent[5..1]
-- Retrieval info: USED_PORT: done 0 0 0 0 OUTPUT NODEFVAL done
-- Retrieval info: USED_PORT: writeenable 0 0 0 0 OUTPUT NODEFVAL writeenable
-- Retrieval info: USED_PORT: direction 0 0 0 0 OUTPUT NODEFVAL direction
-- Retrieval info: CONNECT: @sysclk 0 0 0 0 sysclk 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @go 0 0 0 0 go 0 0 0 0
-- Retrieval info: CONNECT: done 0 0 0 0 @done 0 0 0 0
-- Retrieval info: CONNECT: @realdatain 0 0 16 1 realdatain 0 0 16 1
-- Retrieval info: CONNECT: @imagdatain 0 0 16 1 imagdatain 0 0 16 1
-- Retrieval info: CONNECT: realdataout 0 0 16 1 @realdataout 0 0 16 1
-- Retrieval info: CONNECT: imagdataout 0 0 16 1 @imagdataout 0 0 16 1
-- Retrieval info: CONNECT: @realtwid 0 0 16 1 realtwid 0 0 16 1
-- Retrieval info: CONNECT: @imagtwid 0 0 16 1 imagtwid 0 0 16 1
-- Retrieval info: CONNECT: exponent 0 0 5 1 @exponent 0 0 5 1
-- Retrieval info: CONNECT: readaddress 0 0 8 1 @readaddress 0 0 8 1
-- Retrieval info: CONNECT: writeaddress 0 0 8 1 @writeaddress 0 0 8 1
-- Retrieval info: CONNECT: twidaddress 0 0 8 1 @twidaddress 0 0 8 1
-- Retrieval info: CONNECT: writeenable 0 0 0 0 @writeenable 0 0 0 0
-- Retrieval info: CONNECT: direction 0 0 0 0 @direction 0 0 0 0
